`timescale 1ns / 1ps
module memory(Address, Data);
    input [3:0]Address;
    output [127:0]Data;
    reg [127:0] mem [0:15];
    
    initial 
	begin
		mem[0]  = 128'h54776F204F6E65204E696E652054776F;
		mem[1]  = 128'h03610938AACE8EA1F749B765EEAD464F;
		mem[2]  = 128'hC377E35A37B1BE9D74C5B166769B2F5A;
		mem[3]  = 128'hF5C3C0C5DD4ADE302FA3AFD2E68B09F0;
		mem[4]  = 128'hAD3505D474AA1052A26CC4E51C272B5B;
		mem[5]  = 128'h195C6F2AED81727999B32B9401ECB6E9;
		mem[6]  = 128'hBBC0B840965AE54BB36E227186F81307;
		mem[7]  = 128'h7854B8891BDF022BC28C3BC17F7C50B5;
		mem[8]  = 128'hB5DB295C6EEAC5BF7724767F5E01F2A0;
		mem[9]  = 128'h9F231CAD332DCDDCBD8D7E091F24CB36;
		mem[10] = 128'h1D6DBBABCFB7988D8EF912F76883CDC1;
		mem[11] = 128'h999A215B60A382880D4D9EE16CBB9F52;
		mem[12] = 128'h583F61F14546D1E88A8E1E3A1AD67339;
		mem[13] = 128'hC0BD6F85026FD679EA339E8119B721D3;
		mem[14] = 128'h59BF9E2822DB7B53C839D1D185486D36;
		mem[15] = 128'hD96421AF4B1A50E869E80612A84FCED3;
    end
   
    assign Data = mem[Address][127:0];

endmodule   