`timescale 1ns / 1ps

// just a giant case statement
module sub_byte(SUB_ADDR, SUB_BYTE);
    input [7:0] SUB_ADDR;
    output reg [7:0] SUB_BYTE;
    always @(SUB_ADDR) begin
        case(SUB_ADDR)
            0: SUB_BYTE = 8'h63;
            1: SUB_BYTE = 8'h7c;
            2: SUB_BYTE = 8'h77;
            3: SUB_BYTE = 8'h7b;
            4: SUB_BYTE = 8'hf2;
            5: SUB_BYTE = 8'h6b;
            6: SUB_BYTE = 8'h6f;
            7: SUB_BYTE = 8'hc5;
            8: SUB_BYTE = 8'h30;
            9: SUB_BYTE = 8'h01;
            10: SUB_BYTE = 8'h67;
            11: SUB_BYTE = 8'h2b;
            12: SUB_BYTE = 8'hfe;
            13: SUB_BYTE = 8'hd7;
            14: SUB_BYTE = 8'hab;
            15: SUB_BYTE = 8'h76;
            16: SUB_BYTE = 8'hca;
            17: SUB_BYTE = 8'h82;
            18: SUB_BYTE = 8'hc9;
            19: SUB_BYTE = 8'h7d;
            20: SUB_BYTE = 8'hfa;
            21: SUB_BYTE = 8'h59;
            22: SUB_BYTE = 8'h47;
            23: SUB_BYTE = 8'hf0;
            24: SUB_BYTE = 8'had;
            25: SUB_BYTE = 8'hd4;
            26: SUB_BYTE = 8'ha2;
            27: SUB_BYTE = 8'haf;
            28: SUB_BYTE = 8'h9c;
            29: SUB_BYTE = 8'ha4;
            30: SUB_BYTE = 8'h72;
            31: SUB_BYTE = 8'hc0;
            32: SUB_BYTE = 8'hb7;
            33: SUB_BYTE = 8'hfd;
            34: SUB_BYTE = 8'h93;
            35: SUB_BYTE = 8'h26;
            36: SUB_BYTE = 8'h36;
            37: SUB_BYTE = 8'h3f;
            38: SUB_BYTE = 8'hf7;
            39: SUB_BYTE = 8'hcc;
            40: SUB_BYTE = 8'h34;
            41: SUB_BYTE = 8'ha5;
            42: SUB_BYTE = 8'he5;
            43: SUB_BYTE = 8'hf1;
            44: SUB_BYTE = 8'h71;
            45: SUB_BYTE = 8'hd8;
            46: SUB_BYTE = 8'h31;
            47: SUB_BYTE = 8'h15;
            48: SUB_BYTE = 8'h04;
            49: SUB_BYTE = 8'hc7;
            50: SUB_BYTE = 8'h23;
            51: SUB_BYTE = 8'hc3;
            52: SUB_BYTE = 8'h18;
            53: SUB_BYTE = 8'h96;
            54: SUB_BYTE = 8'h05;
            55: SUB_BYTE = 8'h9a;
            56: SUB_BYTE = 8'h07;
            57: SUB_BYTE = 8'h12;
            58: SUB_BYTE = 8'h80;
            59: SUB_BYTE = 8'he2;
            60: SUB_BYTE = 8'heb;
            61: SUB_BYTE = 8'h27;
            62: SUB_BYTE = 8'hb2;
            63: SUB_BYTE = 8'h75;
            64: SUB_BYTE = 8'h09;
            65: SUB_BYTE = 8'h83;
            66: SUB_BYTE = 8'h2c;
            67: SUB_BYTE = 8'h1a;
            68: SUB_BYTE = 8'h1b;
            69: SUB_BYTE = 8'h6e;
            70: SUB_BYTE = 8'h5a;
            71: SUB_BYTE = 8'ha0;
            72: SUB_BYTE = 8'h52;
            73: SUB_BYTE = 8'h3b;
            74: SUB_BYTE = 8'hd6;
            75: SUB_BYTE = 8'hb3;
            76: SUB_BYTE = 8'h29;
            77: SUB_BYTE = 8'he3;
            78: SUB_BYTE = 8'h2f;
            79: SUB_BYTE = 8'h84;
            80: SUB_BYTE = 8'h53;
            81: SUB_BYTE = 8'hd1;
            82: SUB_BYTE = 8'h00;
            83: SUB_BYTE = 8'hed;
            84: SUB_BYTE = 8'h20;
            85: SUB_BYTE = 8'hfc;
            86: SUB_BYTE = 8'hb1;
            87: SUB_BYTE = 8'h5b;
            88: SUB_BYTE = 8'h6a;
            89: SUB_BYTE = 8'hcb;
            90: SUB_BYTE = 8'hbe;
            91: SUB_BYTE = 8'h39;
            92: SUB_BYTE = 8'h4a;
            93: SUB_BYTE = 8'h4c;
            94: SUB_BYTE = 8'h58;
            95: SUB_BYTE = 8'hcf;
            96: SUB_BYTE = 8'hd0;
            97: SUB_BYTE = 8'hef;
            98: SUB_BYTE = 8'haa;
            99: SUB_BYTE = 8'hfb;
            100: SUB_BYTE = 8'h43;
            101: SUB_BYTE = 8'h4d;
            102: SUB_BYTE = 8'h33;
            103: SUB_BYTE = 8'h85;
            104: SUB_BYTE = 8'h45;
            105: SUB_BYTE = 8'hf9;
            106: SUB_BYTE = 8'h02;
            107: SUB_BYTE = 8'h7f;
            108: SUB_BYTE = 8'h50;
            109: SUB_BYTE = 8'h3c;
            110: SUB_BYTE = 8'h9f;
            111: SUB_BYTE = 8'ha8;
            112: SUB_BYTE = 8'h51;
            113: SUB_BYTE = 8'ha3;
            114: SUB_BYTE = 8'h40;
            115: SUB_BYTE = 8'h8f;
            116: SUB_BYTE = 8'h92;
            117: SUB_BYTE = 8'h9d;
            118: SUB_BYTE = 8'h38;
            119: SUB_BYTE = 8'hf5;
            120: SUB_BYTE = 8'hbc;
            121: SUB_BYTE = 8'hb6;
            122: SUB_BYTE = 8'hda;
            123: SUB_BYTE = 8'h21;
            124: SUB_BYTE = 8'h10;
            125: SUB_BYTE = 8'hff;
            126: SUB_BYTE = 8'hf3;
            127: SUB_BYTE = 8'hd2;
            128: SUB_BYTE = 8'hcd;
            129: SUB_BYTE = 8'h0c;
            130: SUB_BYTE = 8'h13;
            131: SUB_BYTE = 8'hec;
            132: SUB_BYTE = 8'h5f;
            133: SUB_BYTE = 8'h97;
            134: SUB_BYTE = 8'h44;
            135: SUB_BYTE = 8'h17;
            136: SUB_BYTE = 8'hc4;
            137: SUB_BYTE = 8'ha7;
            138: SUB_BYTE = 8'h7e;
            139: SUB_BYTE = 8'h3d;
            140: SUB_BYTE = 8'h64;
            141: SUB_BYTE = 8'h5d;
            142: SUB_BYTE = 8'h19;
            143: SUB_BYTE = 8'h73;
            144: SUB_BYTE = 8'h60;
            145: SUB_BYTE = 8'h81;
            146: SUB_BYTE = 8'h4f;
            147: SUB_BYTE = 8'hdc;
            148: SUB_BYTE = 8'h22;
            149: SUB_BYTE = 8'h2a;
            150: SUB_BYTE = 8'h90;
            151: SUB_BYTE = 8'h88;
            152: SUB_BYTE = 8'h46;
            153: SUB_BYTE = 8'hee;
            154: SUB_BYTE = 8'hb8;
            155: SUB_BYTE = 8'h14;
            156: SUB_BYTE = 8'hde;
            157: SUB_BYTE = 8'h5e;
            158: SUB_BYTE = 8'h0b;
            159: SUB_BYTE = 8'hdb;
            160: SUB_BYTE = 8'he0;
            161: SUB_BYTE = 8'h32;
            162: SUB_BYTE = 8'h3a;
            163: SUB_BYTE = 8'h0a;
            164: SUB_BYTE = 8'h49;
            165: SUB_BYTE = 8'h06;
            166: SUB_BYTE = 8'h24;
            167: SUB_BYTE = 8'h5c;
            168: SUB_BYTE = 8'hc2;
            169: SUB_BYTE = 8'hd3;
            170: SUB_BYTE = 8'hac;
            171: SUB_BYTE = 8'h62;
            172: SUB_BYTE = 8'h91;
            173: SUB_BYTE = 8'h95;
            174: SUB_BYTE = 8'he4;
            175: SUB_BYTE = 8'h79;
            176: SUB_BYTE = 8'he7;
            177: SUB_BYTE = 8'hc8;
            178: SUB_BYTE = 8'h37;
            179: SUB_BYTE = 8'h6d;
            180: SUB_BYTE = 8'h8d;
            181: SUB_BYTE = 8'hd5;
            182: SUB_BYTE = 8'h4e;
            183: SUB_BYTE = 8'ha9;
            184: SUB_BYTE = 8'h6c;
            185: SUB_BYTE = 8'h56;
            186: SUB_BYTE = 8'hf4;
            187: SUB_BYTE = 8'hea;
            188: SUB_BYTE = 8'h65;
            189: SUB_BYTE = 8'h7a;
            190: SUB_BYTE = 8'hae;
            191: SUB_BYTE = 8'h08;
            192: SUB_BYTE = 8'hba;
            193: SUB_BYTE = 8'h78;
            194: SUB_BYTE = 8'h25;
            195: SUB_BYTE = 8'h2e;
            196: SUB_BYTE = 8'h1c;
            197: SUB_BYTE = 8'ha6;
            198: SUB_BYTE = 8'hb4;
            199: SUB_BYTE = 8'hc6;
            200: SUB_BYTE = 8'he8;
            201: SUB_BYTE = 8'hdd;
            202: SUB_BYTE = 8'h74;
            203: SUB_BYTE = 8'h1f;
            204: SUB_BYTE = 8'h4b;
            205: SUB_BYTE = 8'hbd;
            206: SUB_BYTE = 8'h8b;
            207: SUB_BYTE = 8'h8a;
            208: SUB_BYTE = 8'h70;
            209: SUB_BYTE = 8'h3e;
            210: SUB_BYTE = 8'hb5;
            211: SUB_BYTE = 8'h66;
            212: SUB_BYTE = 8'h48;
            213: SUB_BYTE = 8'h03;
            214: SUB_BYTE = 8'hf6;
            215: SUB_BYTE = 8'h0e;
            216: SUB_BYTE = 8'h61;
            217: SUB_BYTE = 8'h35;
            218: SUB_BYTE = 8'h57;
            219: SUB_BYTE = 8'hb9;
            220: SUB_BYTE = 8'h86;
            221: SUB_BYTE = 8'hc1;
            222: SUB_BYTE = 8'h1d;
            223: SUB_BYTE = 8'h9e;
            224: SUB_BYTE = 8'he1;
            225: SUB_BYTE = 8'hf8;
            226: SUB_BYTE = 8'h98;
            227: SUB_BYTE = 8'h11;
            228: SUB_BYTE = 8'h69;
            229: SUB_BYTE = 8'hd9;
            230: SUB_BYTE = 8'h8e;
            231: SUB_BYTE = 8'h94;
            232: SUB_BYTE = 8'h9b;
            233: SUB_BYTE = 8'h1e;
            234: SUB_BYTE = 8'h87;
            235: SUB_BYTE = 8'he9;
            236: SUB_BYTE = 8'hce;
            237: SUB_BYTE = 8'h55;
            238: SUB_BYTE = 8'h28;
            239: SUB_BYTE = 8'hdf;
            240: SUB_BYTE = 8'h8c;
            241: SUB_BYTE = 8'ha1;
            242: SUB_BYTE = 8'h89;
            243: SUB_BYTE = 8'h0d;
            244: SUB_BYTE = 8'hbf;
            245: SUB_BYTE = 8'he6;
            246: SUB_BYTE = 8'h42;
            247: SUB_BYTE = 8'h68;
            248: SUB_BYTE = 8'h41;
            249: SUB_BYTE = 8'h99;
            250: SUB_BYTE = 8'h2d;
            251: SUB_BYTE = 8'h0f;
            252: SUB_BYTE = 8'hb0;
            253: SUB_BYTE = 8'h54;
            254: SUB_BYTE = 8'hbb;
            255: SUB_BYTE = 8'h16;
       endcase
   end
endmodule
